`default_nettype none

module top_module(
    input clk
);



endmodule